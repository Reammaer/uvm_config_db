

package uvm_class_pkg;

    `include "uvm_macros.svh"
    import uvm_pkg::*;

    `include "uvm_classes/agent.sv"
    `include "uvm_classes/environment.sv"
    `include "uvm_classes/base_test.sv"

endpackage: uvm_class_pkg